`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Project Name: RoadRash
// Engineer: Venkata Hemanth Tulimilli
// 
// Create Date: 05/01/2015 01:37:55 AM
// Module Name: icon_module
// Target Devices: Nexys4DDR
// Description: This module takes the input from main controller and then display respective icons depending on those inputs.
// This module is made to display 5 layers with 16 icons in total each depending on the control inputs generated by an LFSR 
// or any other random number generator logic. 
// 5 layers are background layer, bike display layer, two car icon layers, score layer, and speed layer.
// each and every icon displaying logic is implemented in parallel using different always blocks
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// This file is totally dependent on main logic file where we gives out control signals.
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module icon_module (
        input sysreset,
        input sysclk,
        input [9:0]	 bike_col_position,
        input [9:0]  left_car_row, left_car_column, right_car_row, right_car_column, middle_car_row, middle_car_column,
        input [2:0]  left_car_icon_num_port, right_car_icon_num_port, middle_car_icon_num_port, background_num,
        input [10:0] pixel_row,
        input [10:0] pixel_column,
        input [3:0] speed_hunds,
        input [3:0] speed_tens,
        input [3:0] speed_ones,
        input [3:0] score_ones,
        input [3:0] score_tens,
        input [3:0] score_hunds,
        input [3:0] score_thous,
        input [3:0] score_tenthous,
        input [3:0] score_hundthous,

        output reg [7:0] icon,
        output reg       collision_flag,
        output reg [15:0] leds
    );
    
    // local parameters for bike icon on the background
    localparam  BIKE_ROW_START      = 10'd485;
    localparam  BIKE_ROW_END        = 10'd741;
    localparam  BIKE_COL_PIXELS     = 10'd116;
    localparam  BIKE_COL_CHANGE     = 10'd8;
    
    // local parameters for icon sizes for different car sizes to implement 3D illusion
    localparam      ICON_NUM_1          = 10'd16;
    localparam      ICON_NUM_2          = 10'd32;
    localparam      ICON_NUM_3          = 10'd64;
    localparam      ICON_NUM_4          = 10'd128;
    localparam      ICON_NUM_5          = 10'd256;
    
	// score icon and 6 score digits icon row and column start and end pixel values
    localparam      SCORE_ROW_START         = 10'd16;
    localparam      SCORE_COL_START         = 10'd418;
    localparam      SCORE_ROW_END           = 10'd31;
    localparam      SCORE_COL_END           = 10'd481;
    localparam      SCORE_NUM1_ROW_START    = 10'd16;
    localparam      SCORE_NUM1_COL_START    = 10'd490;
    localparam      SCORE_NUM1_ROW_END      = 10'd31;
    localparam      SCORE_NUM1_COL_END      = 10'd505;
    localparam      SCORE_NUM2_ROW_START    = 10'd16;
    localparam      SCORE_NUM2_COL_START    = 10'd510;
    localparam      SCORE_NUM2_ROW_END      = 10'd31;
    localparam      SCORE_NUM2_COL_END      = 10'd525;
    localparam      SCORE_NUM3_ROW_START    = 10'd16;
    localparam      SCORE_NUM3_COL_START    = 10'd530;
    localparam      SCORE_NUM3_ROW_END      = 10'd31;
    localparam      SCORE_NUM3_COL_END      = 10'd545;
    localparam      SCORE_NUM4_ROW_START    = 10'd16;
    localparam      SCORE_NUM4_COL_START    = 10'd550;
    localparam      SCORE_NUM4_ROW_END      = 10'd31;
    localparam      SCORE_NUM4_COL_END      = 10'd565;
    localparam      SCORE_NUM5_ROW_START    = 10'd16;
    localparam      SCORE_NUM5_COL_START    = 10'd570;
    localparam      SCORE_NUM5_ROW_END      = 10'd31;
    localparam      SCORE_NUM5_COL_END      = 10'd585;
    localparam      SCORE_NUM6_ROW_START    = 10'd16;
    localparam      SCORE_NUM6_COL_START    = 10'd590;
    localparam      SCORE_NUM6_ROW_END      = 10'd31;
    localparam      SCORE_NUM6_COL_END      = 10'd605;
    
	// speed icon, numbers and MPH icon row and column start and end pixel values
    localparam      SPEED_ROW_START         = 10'd48;
    localparam      SPEED_COL_START         = 10'd428;
    localparam      SPEED_ROW_END           = 10'd63;
    localparam      SPEED_COL_END           = 10'd491;
    localparam      SPEED_NUM1_ROW_START    = 10'd48;
    localparam      SPEED_NUM1_COL_START    = 10'd500;
    localparam      SPEED_NUM1_ROW_END      = 10'd63;
    localparam      SPEED_NUM1_COL_END      = 10'd515;
    localparam      SPEED_NUM2_ROW_START    = 10'd48;
    localparam      SPEED_NUM2_COL_START    = 10'd520;
    localparam      SPEED_NUM2_ROW_END      = 10'd63;
    localparam      SPEED_NUM2_COL_END      = 10'd535;
    localparam      SPEED_NUM3_ROW_START    = 10'd48;
    localparam      SPEED_NUM3_COL_START    = 10'd540;
    localparam      SPEED_NUM3_ROW_END      = 10'd63;
    localparam      SPEED_NUM3_COL_END      = 10'd555;
    localparam      MPH_ROW_START           = 10'd48;
    localparam      MPH_COL_START           = 10'd564;
    localparam      MPH_ROW_END             = 10'd63;
    localparam      MPH_COL_END             = 10'd595;

	// Local declarations both wire and registers of different lengths
    wire [9:0] LocX, LocY, BotInfo;
    wire reset;
    wire [7:0]  background1_value_wire, background2_value_wire, background3_value_wire, background4_value_wire,
                background5_value_wire, background6_value_wire, background7_value_wire, background8_value_wire;
    wire [7:0] gameover_value_wire;
    wire [7:0] bike_value;
    reg [7:0] left_car_value, middle_car_value, right_car_value, dout3;
    reg [7:0] background_value;
    wire clk;
	reg [15:0] background_addr;
	reg [13:0] gameover_addr;
	reg [14:0] bike_addr;
	reg [9:0] speed_addr;
	reg [9:0] score_addr;
	reg [7:0] number_addr;
	reg [8:0] mph_addr;
	
	reg [7:0] num0_addr;
	wire [7:0] num0_value_wire;
    reg [7:0] num0_value;
    assign num0_value_wire = num0_value;
	
	reg [7:0] num1_addr;
	wire [7:0] num1_value_wire;
    reg [7:0] num1_value;
    assign num1_value_wire = num1_value;
	
	reg [7:0] num2_addr;
	wire [7:0] num2_value_wire;
    reg [7:0] num2_value;
    assign num2_value_wire = num2_value;
	
	reg [7:0] num3_addr;
	wire [7:0] num3_value_wire;
    reg [7:0] num3_value;
    assign num3_value_wire = num3_value;
	
	reg [7:0] num4_addr;
	wire [7:0] num4_value_wire;
    reg [7:0] num4_value;
    assign num4_value_wire = num4_value;
	
	reg [7:0] num5_addr;
	wire [7:0] num5_value_wire;
    reg [7:0] num5_value;
    assign num5_value_wire = num5_value;
	
	reg [7:0] num6_addr;
	wire [7:0] num6_value_wire;
    reg [7:0] num6_value;
    assign num6_value_wire = num6_value;
	
	reg [7:0] num7_addr;
	wire [7:0] num7_value_wire;
    reg [7:0] num7_value;
    assign num7_value_wire = num7_value;
	
	reg [7:0] num8_addr;
	wire [7:0] num8_value_wire;
    reg [7:0] num8_value;
    assign num8_value_wire = num8_value;
	
	reg [7:0] num9_addr;
	wire [7:0] num9_value_wire;
	reg [7:0] num9_value;
    assign num9_value_wire = num9_value;
	
	reg [15:0] left_car5_addr, middle_car5_addr, right_car5_addr;
    reg [13:0] left_car4_addr, middle_car4_addr, right_car4_addr;
    reg [11:0] left_car3_addr, middle_car3_addr, right_car3_addr;
    reg [9:0] left_car2_addr, middle_car2_addr, right_car2_addr;
    reg [7:0] left_car1_addr, middle_car1_addr, right_car1_addr;

    wire [2:0]  left_car_icon_num, right_car_icon_num, middle_car_icon_num;
    assign left_car_icon_num = left_car_icon_num_port;
    assign right_car_icon_num = right_car_icon_num_port;
    assign middle_car_icon_num = middle_car_icon_num_port;
    
    wire [7:0] left_car1_value_wire, left_car2_value_wire, left_car3_value_wire, left_car4_value_wire, left_car5_value_wire;
    wire [7:0] middle_car1_value_wire, middle_car2_value_wire, middle_car3_value_wire, middle_car4_value_wire, middle_car5_value_wire;
    wire [7:0] right_car1_value_wire, right_car2_value_wire, right_car3_value_wire, right_car4_value_wire, right_car5_value_wire;
    wire [7:0] speed_value_wire, score_value_wire, number_value_wire, mph_value_wire;
    reg [7:0]   background1_value, background2_value, background3_value, background4_value, 
                background5_value, background6_value, background7_value, background8_value;
    reg [7:0] gameover_value;
    reg [7:0] speed_value, score_value, mph_value,
              score_num1_value,
              score_num2_value,
              score_num3_value,
              score_num4_value,
              score_num5_value,
              score_num6_value,
              speed_num1_value,
              speed_num2_value,
              speed_num3_value;
    
	reg [7:0] left_car5_value, middle_car5_value, right_car5_value;
    reg [7:0] left_car4_value, middle_car4_value, right_car4_value;
    reg [7:0] left_car3_value, middle_car3_value, right_car3_value;
    reg [7:0] left_car2_value, middle_car2_value, right_car2_value;
    reg [7:0] left_car1_value, middle_car1_value, right_car1_value;
	reg [7:0]  temp_bike_row_addr;
	reg [6:0]  temp_bike_col_addr;
	reg [9:0]  temp_left_car_row_addr, temp_left_car_col_addr,
	           temp_left_car1_row_addr, temp_left_car1_col_addr,
	           temp_left_car2_row_addr, temp_left_car2_col_addr,
	           temp_left_car3_row_addr, temp_left_car3_col_addr,
	           temp_left_car4_row_addr, temp_left_car4_col_addr,
	           temp_left_car5_row_addr, temp_left_car5_col_addr;
	reg [9:0]  temp_middle_car_row_addr, temp_middle_car_col_addr,
	           temp_middle_car1_row_addr, temp_middle_car1_col_addr,
	           temp_middle_car2_row_addr, temp_middle_car2_col_addr,
	           temp_middle_car3_row_addr, temp_middle_car3_col_addr,
	           temp_middle_car4_row_addr, temp_middle_car4_col_addr,
	           temp_middle_car5_row_addr, temp_middle_car5_col_addr;
	reg [9:0]  temp_right_car_row_addr, temp_right_car_col_addr,
	           temp_right_car1_row_addr, temp_right_car1_col_addr,
	           temp_right_car2_row_addr, temp_right_car2_col_addr,
	           temp_right_car3_row_addr, temp_right_car3_col_addr,
	           temp_right_car4_row_addr, temp_right_car4_col_addr,
	           temp_right_car5_row_addr, temp_right_car5_col_addr;
	reg [9:0]  temp_speed_num_row_addr, temp_speed_num_col_addr,
	           temp_score_num_row_addr, temp_score_num_col_addr,
	           temp_speed_row_addr, temp_speed_col_addr,
               temp_score_row_addr, temp_score_col_addr,
               temp_mph_row_addr, temp_mph_col_addr;
	reg        bike_flag;
    reg        left_car_display_flag, 
			   right_car_display_flag, 
			   middle_car_display_flag, 
			   score_display_flag, 
			   speed_display_flag, 
			   mph_display_flag,
               score_num1_display_flag,
               score_num2_display_flag,
               score_num3_display_flag,
               score_num4_display_flag,
               score_num5_display_flag,
               score_num6_display_flag,
               speed_num1_display_flag,
               speed_num2_display_flag,
               speed_num3_display_flag;
    
    assign speed_value_wire = speed_value;
    assign score_value_wire = score_value;
    assign num0_value_wire = num0_value;
    assign num1_value_wire = num1_value;
    assign num2_value_wire = num2_value;
    assign num3_value_wire = num3_value;
    assign num4_value_wire = num4_value;
    assign num5_value_wire = num5_value;
    assign num6_value_wire = num6_value;
    assign num7_value_wire = num7_value;
    assign num8_value_wire = num8_value;
    assign num9_value_wire = num9_value;
    assign mph_value_wire = mph_value;
    
    assign reset = sysreset;
    assign clk = sysclk;
    assign left_car1_value_wire = left_car1_value;
    assign left_car2_value_wire = left_car2_value;
    assign left_car3_value_wire = left_car3_value;
    assign left_car4_value_wire = left_car4_value;
    assign left_car5_value_wire = left_car5_value;

    assign middle_car1_value_wire = middle_car1_value;
    assign middle_car2_value_wire = middle_car2_value;
    assign middle_car3_value_wire = middle_car3_value;
    assign middle_car4_value_wire = middle_car4_value;
    assign middle_car5_value_wire = middle_car5_value;

    assign right_car1_value_wire = right_car1_value;
    assign right_car2_value_wire = right_car2_value;
    assign right_car3_value_wire = right_car3_value;
    assign right_car4_value_wire = right_car4_value;
    assign right_car5_value_wire = right_car5_value;
    
    assign background1_value_wire = background1_value;
    assign background2_value_wire = background2_value;
    assign background3_value_wire = background3_value;
    assign background4_value_wire = background4_value;
    assign background5_value_wire = background5_value;
    assign background6_value_wire = background6_value;
    assign background7_value_wire = background7_value;
    assign background8_value_wire = background8_value;
    
    assign gameover_value_wire = gameover_value;

	// ROMs declarations for different images which are to be displayed on the screen
	background1 BACKGROUND1 (
							.clka(clk),
							.addra(background_addr),
							.douta(background1_value_wire)
							); 
    background2 BACKGROUND2 (
							.clka(clk),
							.addra(background_addr),
							.douta(background2_value_wire)
							); 
    background3 BACKGROUND3 (
							.clka(clk),
							.addra(background_addr),
							.douta(background3_value_wire)
							); 
    background4 BACKGROUND4 (
							.clka(clk),
							.addra(background_addr),
							.douta(background4_value_wire)
							); 
	background5 BACKGROUND5 (
							.clka(clk),
							.addra(background_addr),
							.douta(background5_value_wire)
							); 
	background6 BACKGROUND6 (
							.clka(clk),
							.addra(background_addr),
							.douta(background6_value_wire)
							); 
	background7 BACKGROUND7 (
							.clka(clk),
							.addra(background_addr),
							.douta(background7_value_wire)
							); 
	background8 BACKGROUND8 (
							.clka(clk),
							.addra(background_addr),
							.douta(background8_value_wire)
							); 
    score SCORE 			(
							.clka(clk),
							.addra(score_addr),
							.douta(score_value_wire)
							); 
    speed SPEED 			(
							.clka(clk),
							.addra(speed_addr),
							.douta(speed_value_wire)
							); 
    num0 NUM0 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num0_value_wire)
							); 
    num1 NUM1 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num1_value_wire)
							);
    num2 NUM2 				(			
							.clka(clk),
							.addra(number_addr),
							.douta(num2_value_wire)
							); 
    num3 NUM3 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num3_value_wire)
							); 
    num4 NUM4 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num4_value_wire)
							); 
    num5 NUM5 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num5_value_wire)
							); 
    num6 NUM6 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num6_value_wire)
							); 
    num7 NUM7 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num7_value_wire)
							); 
    num8 NUM8 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num8_value_wire)
							); 
    num9 NUM9 				(
							.clka(clk),
							.addra(number_addr),
							.douta(num9_value_wire)
							); 
    mph MPH 				(
							.clka(clk),
							.addra(mph_addr),
							.douta(mph_value_wire)
							); 
	gameover GAMEOVER 		(
							.clka(clk),
							.addra(gameover_addr),
							.douta(gameover_value_wire)
                            ); 
    bike BIKE 				(
							.clka(clk),
							.addra(bike_addr),
							.douta(bike_value)
							); 
    left_car2 LCAR1 		(
							.clka(clk),
							.addra(left_car1_addr),
							.douta(left_car1_value_wire)
							); 
 
    left_car3 LCAR2 		(
							.clka(clk),
							.addra(left_car2_addr),
							.douta(left_car2_value_wire)
							); 
 
    left_car4 LCAR3 		(
							.clka(clk),
							.addra(left_car3_addr),
							.douta(left_car3_value_wire)
							); 
 
    left_car5 LCAR4 		(
							.clka(clk),
							.addra(left_car4_addr),
							.douta(left_car4_value_wire)
							); 
 
    left_car6 LCAR5 		(
							.clka(clk),
							.addra(left_car5_addr),
							.douta(left_car5_value_wire)
							); 
 
    mid_car2 MIDCAR1 		(
							.clka(clk),
							.addra(middle_car1_addr),
							.douta(middle_car1_value_wire)
							); 
 
    mid_car3 MIDCAR2 		(
							.clka(clk),
							.addra(middle_car2_addr),
							.douta(middle_car2_value_wire)
							); 
 
    mid_car4 MIDCAR3 		(
							.clka(clk),
							.addra(middle_car3_addr),
							.douta(middle_car3_value_wire)
							); 
 
    mid_car5 MIDCAR4 		(
							.clka(clk),
							.addra(middle_car4_addr),
							.douta(middle_car4_value_wire)
							); 
 
    mid_car6 MIDCAR5 		(
							.clka(clk),
							.addra(middle_car5_addr),
							.douta(middle_car5_value_wire)
							); 
    right_car2 RIGHTCAR1 	(
                            .clka(clk),
                            .addra(right_car1_addr),
                            .douta(right_car1_value_wire)
                            );
    right_car3 RIGHTCAR2 	(
                            .clka(clk),
                            .addra(right_car2_addr),
                            .douta(right_car2_value_wire)
                            );
    right_car4 RIGHTCAR3 	(
                            .clka(clk),
                            .addra(right_car3_addr),
                            .douta(right_car3_value_wire)
                            );
    right_car5 RIGHTCAR4 	(
                            .clka(clk),
                            .addra(right_car4_addr),
                            .douta(right_car4_value_wire)
                            );
    right_car6 RIGHTCAR5 	(
                            .clka(clk),
                            .addra(right_car5_addr),
                            .douta(right_car5_value_wire)
                            );

//------------------main screen display always block-------------------//
// 
// selecting values to be displayed at each and every pixel based on the flags set in 
// different always blocks written for each and every ICON displays
// hierarchy is defined such that we can see score even if game is over. 
// 
always @(posedge sysclk) begin
    if (reset) begin
        icon <= 8'd0; 
    end
    else if((score_display_flag == 1'b1) && (score_value != 8'd255)) begin
        icon <= score_value;
    end
    else if((score_num1_display_flag == 1'b1) && (score_num1_value != 8'd255)) begin
        icon <= score_num1_value;
    end
    else if((score_num2_display_flag == 1'b1) && (score_num2_value != 8'd255)) begin
        icon <= score_num2_value;
    end
    else if((score_num3_display_flag == 1'b1) && (score_num3_value != 8'd255)) begin
        icon <= score_num3_value;
    end
    else if((score_num4_display_flag == 1'b1) && (score_num4_value != 8'd255)) begin
        icon <= score_num4_value;
    end
    else if((score_num5_display_flag == 1'b1) && (score_num5_value != 8'd255)) begin
        icon <= score_num5_value;
    end
    else if((score_num6_display_flag == 1'b1) && (score_num6_value != 8'd255)) begin
        icon <= score_num6_value;
    end
    else if(collision_flag) begin
        icon <= gameover_value;
    end
    else if((speed_display_flag == 1'b1) && (speed_value != 8'd255)) begin
        icon <= speed_value;
    end
    else if((speed_num1_display_flag == 1'b1) && (speed_num1_value != 8'd255)) begin
        icon <= speed_num1_value;
    end
    else if((speed_num2_display_flag == 1'b1) && (speed_num2_value != 8'd255)) begin
        icon <= speed_num2_value;
    end
    else if((speed_num3_display_flag == 1'b1) && (speed_num3_value != 8'd255)) begin
        icon <= speed_num3_value;
    end
    else if((mph_display_flag == 1'b1) && (mph_value != 8'd255)) begin
        icon <= mph_value;
    end
    else if((left_car_display_flag == 1'b1) && (left_car_value != 8'd255)) begin
        icon <= left_car_value;
    end
    else if((middle_car_display_flag == 1'b1) && (middle_car_value != 8'd255)) begin
        icon <= middle_car_value;
    end
    else if((right_car_display_flag == 1'b1) && (right_car_value != 8'd255)) begin
        icon <= right_car_value;
    end
    else if((bike_flag == 1'b1) && (bike_value != 8'd255)) begin
        icon <= bike_value;
    end
    else begin
        icon <= background_value;
        leds <= 16'hFFFF;
    end
end
     

//------------------speed icon, score icon, mph icon and 10 number icons address select block-------------------//
// 
// calculating addresses for different icons based on pixel position on the screen with 1024x768 resolution
// and enabling corresponding display flags so that those can be displayed in the above always block 
// according to row and column boundaries defined as local parameters in the beginning of file
// 
always @(posedge sysclk) begin
    if (((pixel_row >= SCORE_ROW_START) && (pixel_row <= SCORE_ROW_END)) && ((pixel_column >= SCORE_COL_START) && (pixel_column <= SCORE_COL_END))) begin
        temp_score_col_addr <= pixel_column - SCORE_COL_START;
        temp_score_row_addr <= pixel_row - SCORE_ROW_START;
        score_addr <= {temp_score_row_addr[3:0], temp_score_col_addr[5:0]};
        score_display_flag <= 1'b1;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM1_ROW_START) && (pixel_row <= SCORE_NUM1_ROW_END)) && ((pixel_column >= SCORE_NUM1_COL_START) && (pixel_column <= SCORE_NUM1_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM1_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM1_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b1;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM2_ROW_START) && (pixel_row <= SCORE_NUM2_ROW_END)) && ((pixel_column >= SCORE_NUM2_COL_START) && (pixel_column <= SCORE_NUM2_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM2_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM2_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b1;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM3_ROW_START) && (pixel_row <= SCORE_NUM3_ROW_END)) && ((pixel_column >= SCORE_NUM3_COL_START) && (pixel_column <= SCORE_NUM3_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM3_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM3_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b1;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM4_ROW_START) && (pixel_row <= SCORE_NUM4_ROW_END)) && ((pixel_column >= SCORE_NUM4_COL_START) && (pixel_column <= SCORE_NUM4_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM4_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM4_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b1;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM5_ROW_START) && (pixel_row <= SCORE_NUM5_ROW_END)) && ((pixel_column >= SCORE_NUM5_COL_START) && (pixel_column <= SCORE_NUM5_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM5_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM5_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b1;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SCORE_NUM6_ROW_START) && (pixel_row <= SCORE_NUM6_ROW_END)) && ((pixel_column >= SCORE_NUM6_COL_START) && (pixel_column <= SCORE_NUM6_COL_END))) begin
        temp_score_num_col_addr <= pixel_column - SCORE_NUM6_COL_START;
        temp_score_num_row_addr <= pixel_row - SCORE_NUM6_ROW_START;
        number_addr <= {temp_score_num_row_addr[3:0], temp_score_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b1;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SPEED_ROW_START) && (pixel_row <= SPEED_ROW_END)) && ((pixel_column >= SPEED_COL_START) && (pixel_column <= SPEED_COL_END))) begin
        temp_speed_col_addr <= pixel_column - SPEED_COL_START;
        temp_speed_row_addr <= pixel_row - SPEED_ROW_START;
        speed_addr <= {temp_speed_row_addr[3:0], temp_speed_col_addr[5:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b1;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SPEED_NUM1_ROW_START) && (pixel_row <= SPEED_NUM1_ROW_END)) && ((pixel_column >= SPEED_NUM1_COL_START) && (pixel_column <= SPEED_NUM1_COL_END))) begin
        temp_speed_num_col_addr <= pixel_column - SPEED_NUM1_COL_START;
        temp_speed_num_row_addr <= pixel_row - SPEED_NUM1_ROW_START;
        number_addr <= {temp_speed_num_row_addr[3:0], temp_speed_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b1;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SPEED_NUM2_ROW_START) && (pixel_row <= SPEED_NUM2_ROW_END)) && ((pixel_column >= SPEED_NUM2_COL_START) && (pixel_column <= SPEED_NUM2_COL_END))) begin
        temp_speed_num_col_addr <= pixel_column - SPEED_NUM2_COL_START;
        temp_speed_num_row_addr <= pixel_row - SPEED_NUM2_ROW_START;
        number_addr <= {temp_speed_num_row_addr[3:0], temp_speed_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b1;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= SPEED_NUM3_ROW_START) && (pixel_row <= SPEED_NUM3_ROW_END)) && ((pixel_column >= SPEED_NUM3_COL_START) && (pixel_column <= SPEED_NUM3_COL_END))) begin
        temp_speed_num_col_addr <= pixel_column - SPEED_NUM3_COL_START;
        temp_speed_num_row_addr <= pixel_row - SPEED_NUM3_ROW_START;
        number_addr <= {speed_hunds, temp_speed_num_row_addr[3:0], temp_speed_num_col_addr[3:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b1;
        mph_display_flag <= 1'b0;
    end
    else if (((pixel_row >= MPH_ROW_START) && (pixel_row <= MPH_ROW_END)) && ((pixel_column >= MPH_COL_START) && (pixel_column <= MPH_COL_END))) begin
        temp_mph_col_addr <= pixel_column - MPH_COL_START;
        temp_mph_row_addr <= pixel_row - MPH_ROW_START;
        mph_addr <= {temp_mph_row_addr[3:0], temp_mph_col_addr[4:0]};
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b1;
    end
    else begin
        score_display_flag <= 1'b0;
        speed_display_flag <= 1'b0;
        score_num1_display_flag <= 1'b0;
        score_num2_display_flag <= 1'b0;
        score_num3_display_flag <= 1'b0;
        score_num4_display_flag <= 1'b0;
        score_num5_display_flag <= 1'b0;
        score_num6_display_flag <= 1'b0;
        speed_num1_display_flag <= 1'b0;
        speed_num2_display_flag <= 1'b0;
        speed_num3_display_flag <= 1'b0;
        mph_display_flag <= 1'b0;
    end

end

//------------------speed number1 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "speed_hunds" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       speed_num1_value <= 8'd0;
    end
    else if (speed_hunds == 4'd0) begin
        speed_num1_value <= num0_value;
    end
    else if (speed_hunds == 4'd1) begin
        speed_num1_value <= num1_value;
    end
    else if (speed_hunds == 4'd2) begin
        speed_num1_value <= num2_value;
    end
    else if (speed_hunds == 4'd3) begin
        speed_num1_value <= num3_value;
    end
    else if (speed_hunds == 4'd4) begin
        speed_num1_value <= num4_value;
    end
    else if (speed_hunds == 4'd5) begin
        speed_num1_value <= num5_value;
    end
    else if (speed_hunds == 4'd6) begin
        speed_num1_value <= num6_value;
    end
    else if (speed_hunds == 4'd7) begin
        speed_num1_value <= num7_value;
    end
    else if (speed_hunds == 4'd8) begin
        speed_num1_value <= num8_value;
    end
    else if (speed_hunds == 4'd9) begin
        speed_num1_value <= num9_value;
    end
    else begin
        speed_num1_value <= 8'd255;
    end
end

//------------------speed number2 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "speed_tens" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       speed_num2_value <= 8'd0;
    end
    else if (speed_tens == 4'd0) begin
        speed_num2_value <= num0_value;
    end
    else if (speed_tens == 4'd1) begin
        speed_num2_value <= num1_value;
    end
    else if (speed_tens == 4'd2) begin
        speed_num2_value <= num2_value;
    end
    else if (speed_tens == 4'd3) begin
        speed_num2_value <= num3_value;
    end
    else if (speed_tens == 4'd4) begin
        speed_num2_value <= num4_value;
    end
    else if (speed_tens == 4'd5) begin
        speed_num2_value <= num5_value;
    end
    else if (speed_tens == 4'd6) begin
        speed_num2_value <= num6_value;
    end
    else if (speed_tens == 4'd7) begin
        speed_num2_value <= num7_value;
    end
    else if (speed_tens == 4'd8) begin
        speed_num2_value <= num8_value;
    end
    else if (speed_tens == 4'd9) begin
        speed_num2_value <= num9_value;
    end
    else begin
        speed_num2_value <= 8'd255;
    end
end

//------------------speed number3 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "speed_ones" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       speed_num3_value <= 8'd0;
    end
    else if (speed_ones == 4'd0) begin
        speed_num3_value <= num0_value;
    end
    else if (speed_ones == 4'd1) begin
        speed_num3_value <= num1_value;
    end
    else if (speed_ones == 4'd2) begin
        speed_num3_value <= num2_value;
    end
    else if (speed_ones == 4'd3) begin
        speed_num3_value <= num3_value;
    end
    else if (speed_ones == 4'd4) begin
        speed_num3_value <= num4_value;
    end
    else if (speed_ones == 4'd5) begin
        speed_num3_value <= num5_value;
    end
    else if (speed_ones == 4'd6) begin
        speed_num3_value <= num6_value;
    end
    else if (speed_ones == 4'd7) begin
        speed_num3_value <= num7_value;
    end
    else if (speed_ones == 4'd8) begin
        speed_num3_value <= num8_value;
    end
    else if (speed_ones == 4'd9) begin
        speed_num3_value <= num9_value;
    end
    else begin
        speed_num3_value <= 8'd255;
    end
end

//------------------score number1 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_hundthous" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num1_value <= 8'd0;
    end
    else if (score_hundthous == 4'd0) begin
        score_num1_value <= num0_value;
    end
    else if (score_hundthous == 4'd1) begin
        score_num1_value <= num1_value;
    end
    else if (score_hundthous == 4'd2) begin
        score_num1_value <= num2_value;
    end
    else if (score_hundthous == 4'd3) begin
        score_num1_value <= num3_value;
    end
    else if (score_hundthous == 4'd4) begin
        score_num1_value <= num4_value;
    end
    else if (score_hundthous == 4'd5) begin
        score_num1_value <= num5_value;
    end
    else if (score_hundthous == 4'd6) begin
        score_num1_value <= num6_value;
    end
    else if (score_hundthous == 4'd7) begin
        score_num1_value <= num7_value;
    end
    else if (score_hundthous == 4'd8) begin
        score_num1_value <= num8_value;
    end
    else if (score_hundthous == 4'd9) begin
        score_num1_value <= num9_value;
    end
    else begin
        score_num1_value <= 8'd255;
    end
end

//------------------score number2 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_tenthous" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num2_value <= 8'd0;
    end
    else if (score_tenthous == 4'd0) begin
        score_num2_value <= num0_value;
    end
    else if (score_tenthous == 4'd1) begin
        score_num2_value <= num1_value;
    end
    else if (score_tenthous == 4'd2) begin
        score_num2_value <= num2_value;
    end
    else if (score_tenthous == 4'd3) begin
        score_num2_value <= num3_value;
    end
    else if (score_tenthous == 4'd4) begin
        score_num2_value <= num4_value;
    end
    else if (score_tenthous == 4'd5) begin
        score_num2_value <= num5_value;
    end
    else if (score_tenthous == 4'd6) begin
        score_num2_value <= num6_value;
    end
    else if (score_tenthous == 4'd7) begin
        score_num2_value <= num7_value;
    end
    else if (score_tenthous == 4'd8) begin
        score_num2_value <= num8_value;
    end
    else if (score_tenthous == 4'd9) begin
        score_num2_value <= num9_value;
    end
    else begin
        score_num2_value <= 8'd255;
    end
end

//------------------score number3 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_thous" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num3_value <= 8'd0;
    end
    else if (score_thous == 4'd0) begin
        score_num3_value <= num0_value;
    end
    else if (score_thous == 4'd1) begin
        score_num3_value <= num1_value;
    end
    else if (score_thous == 4'd2) begin
        score_num3_value <= num2_value;
    end
    else if (score_thous == 4'd3) begin
        score_num3_value <= num3_value;
    end
    else if (score_thous == 4'd4) begin
        score_num3_value <= num4_value;
    end
    else if (score_thous == 4'd5) begin
        score_num3_value <= num5_value;
    end
    else if (score_thous == 4'd6) begin
        score_num3_value <= num6_value;
    end
    else if (score_thous == 4'd7) begin
        score_num3_value <= num7_value;
    end
    else if (score_thous == 4'd8) begin
        score_num3_value <= num8_value;
    end
    else if (score_thous == 4'd9) begin
        score_num3_value <= num9_value;
    end
    else begin
        score_num3_value <= 8'd255;
    end
end

//------------------score number4 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_hunds" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num4_value <= 8'd0;
    end
    else if (score_hunds == 4'd0) begin
        score_num4_value <= num0_value;
    end
    else if (score_hunds == 4'd1) begin
        score_num4_value <= num1_value;
    end
    else if (score_hunds == 4'd2) begin
        score_num4_value <= num2_value;
    end
    else if (score_hunds == 4'd3) begin
        score_num4_value <= num3_value;
    end
    else if (score_hunds == 4'd4) begin
        score_num4_value <= num4_value;
    end
    else if (score_hunds == 4'd5) begin
        score_num4_value <= num5_value;
    end
    else if (score_hunds == 4'd6) begin
        score_num4_value <= num6_value;
    end
    else if (score_hunds == 4'd7) begin
        score_num4_value <= num7_value;
    end
    else if (score_hunds == 4'd8) begin
        score_num4_value <= num8_value;
    end
    else if (score_hunds == 4'd9) begin
        score_num4_value <= num9_value;
    end
    else begin
        score_num4_value <= 8'd255;
    end
end

//------------------score number5 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_tens" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num5_value <= 8'd0;
    end
    else if (score_tens == 4'd0) begin
        score_num5_value <= num0_value;
    end
    else if (score_tens == 4'd1) begin
        score_num5_value <= num1_value;
    end
    else if (score_tens == 4'd2) begin
        score_num5_value <= num2_value;
    end
    else if (score_tens == 4'd3) begin
        score_num5_value <= num3_value;
    end
    else if (score_tens == 4'd4) begin
        score_num5_value <= num4_value;
    end
    else if (score_tens == 4'd5) begin
        score_num5_value <= num5_value;
    end
    else if (score_tens == 4'd6) begin
        score_num5_value <= num6_value;
    end
    else if (score_tens == 4'd7) begin
        score_num5_value <= num7_value;
    end
    else if (score_tens == 4'd8) begin
        score_num5_value <= num8_value;
    end
    else if (score_tens == 4'd9) begin
        score_num5_value <= num9_value;
    end
    else begin
        score_num5_value <= 8'd255;
    end
end

//------------------score number6 icon value select block-------------------//
// 
// selecting 8bit colour value of number icon from different ROMs depending on 
// different "score_ones" value coming from main controller block 
// 
always @(posedge clk) begin
    if(reset) begin
       score_num6_value <= 8'd0;
    end
    else if (score_ones == 4'd0) begin
        score_num6_value <= num0_value;
    end
    else if (score_ones == 4'd1) begin
        score_num6_value <= num1_value;
    end
    else if (score_ones == 4'd2) begin
        score_num6_value <= num2_value;
    end
    else if (score_ones == 4'd3) begin
        score_num6_value <= num3_value;
    end
    else if (score_ones == 4'd4) begin
        score_num6_value <= num4_value;
    end
    else if (score_ones == 4'd5) begin
        score_num6_value <= num5_value;
    end
    else if (score_ones == 4'd6) begin
        score_num6_value <= num6_value;
    end
    else if (score_ones == 4'd7) begin
        score_num6_value <= num7_value;
    end
    else if (score_ones == 4'd8) begin
        score_num6_value <= num8_value;
    end
    else if (score_ones == 4'd9) begin
        score_num6_value <= num9_value;
    end
    else begin
        score_num6_value <= 8'd255;
    end
end

//------------------collision detection block-------------------//
// 
// detecting collision flag so to make sure we detect collision occurred and then stop the game
// based on the collision flag. 
// 
// collision detection is achieved by comparing when bike_flag is HIGH as well as any of the 
// car_display_flag is HIGH after eliminating white values in the icons 
// 
always @(posedge sysclk) begin
    if(reset) begin
        collision_flag <= 1'b0;
    end
    else if (((bike_flag == 1'b1) && (bike_value != 8'd255)) && (((left_car_display_flag == 1'b1) && (left_car_value != 8'd255)) || 
                                                                 ((middle_car_display_flag == 1'b1) && (middle_car_value != 8'd255)) ||
                                                                 ((right_car_display_flag == 1'b1) && (right_car_value != 8'd255)))) begin
        collision_flag <= 1'b1;
    end
    else begin
        collision_flag <= collision_flag;
    end
end
     
//------------------background icon value select block-------------------//
// 
// selecting 8bit colour value of background from different ROMs depending on 
// different background_num or collision_flag values coming from main controller block 
// 
always @(posedge sysclk) begin
    if(reset) begin
        background_value <= 8'd0;
    end
    else if (collision_flag) begin
        background_value <= gameover_value;
    end
    else if (background_num == 3'd0) begin
        background_value <= background1_value;
    end
    else if (background_num == 3'd1) begin
        background_value <= background2_value;
    end
    else if (background_num == 3'd2) begin
        background_value <= background3_value;
    end
    else if (background_num == 3'd3) begin
        background_value <= background4_value;
    end
    else if (background_num == 3'd4) begin
        background_value <= background5_value;
    end
    else if (background_num == 3'd5) begin
        background_value <= background6_value;
    end
    else if (background_num == 3'd6) begin
        background_value <= background7_value;
    end
    else if (background_num == 3'd7) begin
        background_value <= background8_value;
    end
    else begin
       background_value <= background1_value;
    end
end

//------------------left car icon value select block-------------------//
// 
// selecting 8bit colour value of left car from different ROMs depending on 
// different left_car_icon_num values coming from main controller block 
// 
always @(posedge sysclk) begin
    if (reset) begin
        left_car_value <= 8'd0;
    end
    else if ((left_car_icon_num == 3'd1) || (left_car_icon_num == 3'd2)) begin
        left_car_value <= left_car2_value_wire;
    end
    else if (left_car_icon_num == 3'd3) begin
        left_car_value <= left_car3_value_wire;
    end
    else if ((left_car_icon_num == 3'd4) || (left_car_icon_num == 3'd5)) begin
        left_car_value <= left_car5_value_wire;
    end
    else begin
        left_car_value <= 8'd15;
    end
end


//------------------left car icon display block-------------------//
// 
// giving address to left car icon ROMs depending on left_icon_num input which comes 
// from main controller block and enabling left_car_display_flag so that 
// main display block above in different always block displays different icons in different layers
// -----left_car_icon_num----------display pixels--------
// |			1, 2					32 x 32         |
// |			  3						64 x 64         |
// |			4, 5				   256 x 256        |
// ------------------------------------------------------
// 
always @(posedge sysclk)	begin
    
    
    if((left_car_icon_num ==  3'd1) || (left_car_icon_num ==  3'd2)) begin
        if(((pixel_row >= left_car_row) && (pixel_row < (left_car_row + ICON_NUM_2))) && ((pixel_column >= left_car_column) && (pixel_column < (left_car_column + ICON_NUM_2)))) begin
            temp_left_car_col_addr <= pixel_column - left_car_column;
            temp_left_car_row_addr <= pixel_row - left_car_row;
            left_car2_addr <= {temp_left_car_row_addr[4:1], temp_left_car_col_addr[4:1]};
            left_car_display_flag <= 1'b1;
        end
        else begin
            left_car_display_flag <= 1'b0;
        end
    end
    else if(left_car_icon_num ==  3'd3) begin
        if(((pixel_row >= left_car_row) && (pixel_row < (left_car_row + ICON_NUM_3))) && ((pixel_column >= left_car_column) && (pixel_column < (left_car_column + ICON_NUM_3)))) begin
            temp_left_car_col_addr <= pixel_column - left_car_column;
            temp_left_car_row_addr <= pixel_row - left_car_row;
            left_car3_addr <= {temp_left_car_row_addr[5:1], temp_left_car_col_addr[5:1]};
            left_car_display_flag <= 1'b1;
        end
        else begin
            left_car_display_flag <= 1'b0;
        end
    end
    else if((left_car_icon_num ==  3'd4) || (left_car_icon_num ==  3'd5)) begin
        if(((pixel_row >= left_car_row) && (pixel_row < (left_car_row + ICON_NUM_5))) && ((pixel_column >= left_car_column) && (pixel_column < (left_car_column + ICON_NUM_5)))) begin
            temp_left_car_col_addr <= pixel_column - left_car_column;
            temp_left_car_row_addr <= pixel_row - left_car_row;
            left_car5_addr <= {temp_left_car_row_addr[7:1], temp_left_car_col_addr[7:1]};
            left_car_display_flag <= 1'b1;
        end
        else begin
            left_car_display_flag <= 1'b0;
        end
    end
    else begin
        temp_left_car_col_addr <= 7'd0;
        temp_left_car_row_addr <= 7'd0;
        left_car1_addr <= 14'd0;
        left_car_display_flag <= 1'b0;
    end
end

//------------------right car icon value select block-------------------//
// 
// selecting 8bit colour value of right car from different ROMs depending on 
// different right_car_icon_num values coming from main controller block 
// 
always @(posedge sysclk) begin
    if (reset) begin
        right_car_value <= 8'd0;
    end
    else if (right_car_icon_num == 3'd1) begin
        right_car_value <= right_car2_value_wire;
    end
    else if (right_car_icon_num == 3'd2) begin
        right_car_value <= right_car2_value_wire;
    end
    else if (right_car_icon_num == 3'd3) begin
        right_car_value <= right_car3_value_wire;
    end
    else if (right_car_icon_num == 3'd4) begin
        right_car_value <= right_car5_value_wire;
    end
    else if (right_car_icon_num == 3'd5) begin
        right_car_value <= right_car5_value_wire;
    end
    else begin
        right_car_value <= 8'd15;
    end
end

//------------------right car icon display block-------------------//
// 
// giving address to right car icon ROMs depending on right_icon_num input which comes 
// from main controller block and enabling right_car_display_flag so that 
// main display block above in different always block displays different icons in different layers
// -----right_car_icon_num----------display pixels-------
// |			1, 2					32 x 32         |
// |			  3						64 x 64         |
// |			4, 5				   256 x 256        |
// ------------------------------------------------------
// 
always @(posedge sysclk)	begin
    
    
    if((right_car_icon_num ==  3'd1) || (right_car_icon_num ==  3'd2)) begin
        if(((pixel_row >= right_car_row) && (pixel_row < (right_car_row + ICON_NUM_2))) && ((pixel_column >= right_car_column) && (pixel_column < (right_car_column + ICON_NUM_2)))) begin
            temp_right_car_col_addr <= pixel_column - right_car_column;
            temp_right_car_row_addr <= pixel_row - right_car_row;
            right_car2_addr <= {temp_right_car_row_addr[4:1], temp_right_car_col_addr[4:1]};
            right_car_display_flag <= 1'b1;
        end
        else begin
            right_car_display_flag <= 1'b0;
        end
    end
    else if(right_car_icon_num ==  3'd3) begin
        if(((pixel_row >= right_car_row) && (pixel_row < (right_car_row + ICON_NUM_3))) && ((pixel_column >= right_car_column) && (pixel_column < (right_car_column + ICON_NUM_3)))) begin
            temp_right_car_col_addr <= pixel_column - right_car_column;
            temp_right_car_row_addr <= pixel_row - right_car_row;
            right_car3_addr <= {temp_right_car_row_addr[5:1], temp_right_car_col_addr[5:1]};
            right_car_display_flag <= 1'b1;
        end
        else begin
            right_car_display_flag <= 1'b0;
        end
    end
    else if((right_car_icon_num ==  3'd4) || (right_car_icon_num ==  3'd5)) begin
        if(((pixel_row >= right_car_row) && (pixel_row < (right_car_row + ICON_NUM_5))) && ((pixel_column >= right_car_column) && (pixel_column < (right_car_column + ICON_NUM_5)))) begin
            temp_right_car_col_addr <= pixel_column - right_car_column;
            temp_right_car_row_addr <= pixel_row - right_car_row;
            right_car5_addr <= {temp_right_car_row_addr[7:1], temp_right_car_col_addr[7:1]};
            right_car_display_flag <= 1'b1;
        end
        else begin
            right_car_display_flag <= 1'b0;
        end
    end
    else begin
        temp_right_car_col_addr <= 7'd0;
        temp_right_car_row_addr <= 7'd0;
        right_car1_addr <= 14'd0;
        right_car_display_flag <= 1'b0;
    end
end

//------------------middle car icon value select block-------------------//
// 
// selecting 8bit colour value of middle car from different ROMs depending on 
// different middle_car_icon_num values coming from main controller block 
// 
always @(posedge sysclk) begin
    if (reset) begin
        middle_car_value <= 8'd0;
    end
    else if ((middle_car_icon_num == 3'd1) || (middle_car_icon_num == 3'd2)) begin
        middle_car_value <= middle_car2_value_wire;
    end
    else if (middle_car_icon_num == 3'd3) begin
        middle_car_value <= middle_car3_value_wire;
    end
    else if (middle_car_icon_num == 3'd4) begin
        middle_car_value <= middle_car4_value_wire;
    end
    else if (middle_car_icon_num == 3'd5) begin
        middle_car_value <= middle_car5_value_wire;
    end
    else begin
        middle_car_value <= 8'd255;
    end
end

//--------------middle car icon address select block----------------//
// 
// giving address to middle car icon ROMs depending on middle_icon_num input which comes 
// from main controller block and enabling middle_car_display_flag so that 
// main display block above in different always block depending on different flags
// -----middle_car_icon_num----------display pixels-----
// |				1, 2				32 x 32		   |
// |				  3					64 x 64		   |
// |				  4				   128 x 128   	   |
// |				  5				   256 x 256   	   |
// -----------------------------------------------------
// 
always @(posedge sysclk)	begin
    if((middle_car_icon_num ==  3'd1) || (middle_car_icon_num ==  3'd2)) begin
        if(((pixel_row >= middle_car_row) && (pixel_row < (middle_car_row + ICON_NUM_2))) && ((pixel_column >= middle_car_column) && (pixel_column < (middle_car_column + ICON_NUM_2)))) begin
            temp_middle_car_col_addr <= pixel_column - middle_car_column;
            temp_middle_car_row_addr <= pixel_row - middle_car_row;
            middle_car2_addr <= {temp_middle_car_row_addr[4:1], temp_middle_car_col_addr[4:1]};
            middle_car_display_flag <= 1'b1;
        end
        else begin
            middle_car_display_flag <= 1'b0;
        end
    end
    else if(middle_car_icon_num ==  3'd3) begin
        if(((pixel_row >= middle_car_row) && (pixel_row < (middle_car_row + ICON_NUM_3))) && ((pixel_column >= middle_car_column) && (pixel_column < (middle_car_column + ICON_NUM_3)))) begin
            temp_middle_car_col_addr <= pixel_column - middle_car_column;
            temp_middle_car_row_addr <= pixel_row - middle_car_row;
            middle_car3_addr <= {temp_middle_car_row_addr[5:1], temp_middle_car_col_addr[5:1]};
            middle_car_display_flag <= 1'b1;
        end
        else begin
            middle_car_display_flag <= 1'b0;
        end
    end
    else if(middle_car_icon_num ==  3'd4) begin
        if(((pixel_row >= middle_car_row) && (pixel_row < (middle_car_row + ICON_NUM_4))) && ((pixel_column >= middle_car_column) && (pixel_column < (middle_car_column + ICON_NUM_4)))) begin
            temp_middle_car_col_addr <= pixel_column - middle_car_column;
            temp_middle_car_row_addr <= pixel_row - middle_car_row;
            middle_car4_addr <= {temp_middle_car_row_addr[6:1], temp_middle_car_col_addr[6:1]};
            middle_car_display_flag <= 1'b1;
        end
        else begin
            middle_car_display_flag <= 1'b0;
        end
    end
    else if(middle_car_icon_num ==  3'd5) begin
        if(((pixel_row >= middle_car_row) && (pixel_row < (middle_car_row + ICON_NUM_5))) && ((pixel_column >= middle_car_column) && (pixel_column < (middle_car_column + ICON_NUM_5)))) begin
            temp_middle_car_col_addr <= pixel_column - middle_car_column;
            temp_middle_car_row_addr <= pixel_row - middle_car_row;
            middle_car5_addr <= {temp_middle_car_row_addr[7:1], temp_middle_car_col_addr[7:1]};
            middle_car_display_flag <= 1'b1;
        end
        else begin
            middle_car_display_flag <= 1'b0;
        end
    end
    else begin
        temp_middle_car_col_addr <= 7'd0;
        temp_middle_car_row_addr <= 7'd0;
        middle_car1_addr <= 14'd0;
        middle_car_display_flag <= 1'b0;
    end
end

//------------------bike address select block-------------------//
//
// checking the pixels where the bike icon should be displayed
// and enabling bike flag to display on the screen or VGA display
// here always bike row is fixed where as column position is going to
// vary according to logic implemented in main logic controller.
//
always @(posedge sysclk) begin
    if(((pixel_row >= BIKE_ROW_START) && (pixel_row < BIKE_ROW_END)) && ((pixel_column >= bike_col_position) && (pixel_column <( bike_col_position + BIKE_COL_PIXELS)))) begin
        temp_bike_col_addr <= pixel_column - bike_col_position;
        temp_bike_row_addr <= pixel_row - BIKE_ROW_START;
        bike_addr <= {temp_bike_row_addr, temp_bike_col_addr};
        bike_flag <= 1'b1;
    end
    else begin
        temp_bike_col_addr <= 7'd0;
        temp_bike_row_addr <= 8'd0;
        bike_addr <= 15'd0;
        bike_flag <= 1'b0;
    end
end

//------------------background icon display block-------------------//
// 
// giving address to background icons ROMs for both backgrounds 
// as well as game over background image
// 
always @(posedge sysclk) begin
    gameover_addr <= {pixel_row[9:3], pixel_column[9:3]};
    background_addr <= {pixel_row[9:2], pixel_column[9:2]};
end
endmodule